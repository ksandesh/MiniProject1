`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:   
// Design Name: 
// Module Name:    top_level 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module top_level(
    input clk,         // 100mhz clock
    input rst,         // Asynchronous reset, tied to dip switch 0
    output txd,        // RS232 Transmit Data
    input rxd,         // RS232 Recieve Data
    input [1:0] br_cfg, // Baud Rate Configuration, Tied to dip switches 2 and 3
	 output GPIO_LED_0,
	 output GPIO_LED_1,
	 output GPIO_LED_2,
	 output GPIO_LED_3,
	 output GPIO_LED_4,
	 output GPIO_LED_5,
	 output GPIO_LED_6,
	 output GPIO_LED_7
    );
	
	wire iocs;
	wire iorw;
	wire rda;
	wire tbr;
	wire [1:0] ioaddr;
	wire [7:0] databus;
	
	// Instantiate your SPART here
	spart spart0( .clk(clk),
                 .rst(rst),
					  .iocs(iocs),
					  .iorw(iorw),
					  .rda(rda),
					  .tbr(tbr),
					  .ioaddr(ioaddr),
					  .databus(databus),
					  .txd(txd),
					  .rxd(rxd)
					);

	// Instantiate your driver here
	driver driver0( .clk(clk),
	                .rst(rst),
						 .br_cfg(br_cfg),
						 .iocs(iocs),
						 .iorw(iorw),
						 .rda(rda),
						 .tbr(tbr),
						 .ioaddr(ioaddr),
						 .databus(databus),
						 .GPIO_LED_0(GPIO_LED_0),
						 .GPIO_LED_1(GPIO_LED_1),
							.GPIO_LED_2(GPIO_LED_2),
							.GPIO_LED_3(GPIO_LED_3),
							.GPIO_LED_4(GPIO_LED_4),
							.GPIO_LED_5(GPIO_LED_5),
							.GPIO_LED_6(GPIO_LED_6),
							.GPIO_LED_7(GPIO_LED_7)
					 );   
					 
endmodule

